library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity sinus is
  port( rst, h ,amp: std_logic;
    freq : std_logic_vector(3 downto 0);
    mode :std_logic_vector(1 downto 0);
        Vs : out std_logic_vector(9 downto 0) );
end sinus;

architecture rtl of sinus is
  signal sens, signe, eq511, eq0, C1, C2, C3, C4, C5 : std_logic;
  --signal freq : std_logic_vector (3 downto 0);
  signal I : std_logic_vector(8 downto 0);
 --table de valeurs pour g�n�rer un sinus de p�riode 625us
 
  type defsinus is array(0 to 361) of std_logic_vector(8 downto 0);
  constant sinusask :defsinus :=( "000000000", "000000110", "000001011", "000010000", "000010101",
"000011010", "000011111", "000100100", "000101001", "000101110",
"000110011", "000111000", "000111101", "001000010", "001000111",
"001001100", "001010001", "001010110", "001011010", "001011111",
"001100100", "001101001", "001101110", "001110011", "001111000",
"001111101", "010000010", "010000111", "010001011", "010010000",
"010010101", "010011010", "010011111", "010100011", "010101000",
"010101101", "010110010", "010110110", "010111011", "011000000",
"011000100", "011001001", "011001101", "011010010", "011010111",
"011011011", "011100000", "011100100", "011101001", "011101101",
"011110001", "011110110", "011111010", "011111110", "100000011",
"100000111", "100001011", "100010000", "100010100", "100011000",
"100011100", "100100000", "100100100", "100101000", "100101100",
"100110000", "100110100", "100111000", "100111100", "101000000",
"101000100", "101001000", "101001100", "101001111", "101010011",
"101010111", "101011010", "101011110", "101100010", "101100101",
"101101001", "101101100", "101110000", "101110011", "101110110",
"101111010", "101111101", "110000000", "110000011", "110000111",
"110001010", "110001101", "110010000", "110010011", "110010110",
"110011001", "110011100", "110011110", "110100001", "110100100",
"110100111", "110101001", "110101100", "110101111", "110110001",
"110110100", "110110110", "110111000", "110111011", "110111101",
"110111111", "111000010", "111000100", "111000110", "111001000",
"111001010", "111001100", "111001110", "111010000", "111010010",
"111010100", "111010101", "111010111", "111011001", "111011010",
"111011100", "111011110", "111011111", "111100000", "111100010",
"111100011", "111100100", "111100110", "111100111", "111101000",
"111101001", "111101010", "111101011", "111101100", "111101101",
"111101110", "111101111", "111101111", "111110000", "111110001",
"111110001", "111110010", "111110010", "111110011", "111110011",
"111110100", "111110100", "111110100", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );
 
--table de valeurs pour g�n�rer un sinus avec une fr�quence de 697 Hz

constant sinus697 :defsinus :=( "000000000", "000000001", "000000001", "000000001", "000000001",
"000000010", "000000010", "000000010", "000000010", "000000010",
"000000011", "000000011", "000000011", "000000011", "000000100",
"000000100", "000000100", "000000100", "000000100", "000000101",
"000000101", "000000101", "000000101", "000000101", "000000110",
"000000110", "000000110", "000000110", "000000111", "000000111",
"000000111", "000000111", "000000111", "000001000", "000001000",
"000001000", "000001000", "000001001", "000001001", "000001001",
"000001001", "000001001", "000001010", "000001010", "000001010",
"000001010", "000001010", "000001011", "000001011", "000001011",
"000001011", "000001011", "000001100", "000001100", "000001100",
"000001100", "000001101", "000001101", "000001101", "000001101",
"000001101", "000001110", "000001110", "000001110", "000001110",
"000001110", "000001111", "000001111", "000001111", "000001111",
"000001111", "000010000", "000010000", "000010000", "000010000",
"000010001", "000010001", "000010001", "000010001", "000010001",
"000010010", "000010010", "000010010", "000010010", "000010010",
"000010011", "000010011", "000010011", "000010011", "000010011",
"000010100", "000010100", "000010100", "000010100", "000010100",
"000010101", "000010101", "000010101", "000010101", "000010101",
"000010110", "000010110", "000010110", "000010110", "000010110",
"000010111", "000010111", "000010111", "000010111", "000010111",
"000011000", "000011000", "000011000", "000011000", "000011000",
"000011000", "000011001", "000011001", "000011001", "000011001",
"000011001", "000011010", "000011010", "000011010", "000011010",
"000011010", "000011011", "000011011", "000011011", "000011011",
"000011011", "000011011", "000011100", "000011100", "000011100",
"000011100", "000011100", "000011101", "000011101", "000011101",
"000011101", "000011101", "000011101", "000011110", "000011110",
"000011110", "000011110", "000011110", "000011110", "000011111",
"000011111", "000011111", "000011111", "000011111", "000100000",
"000100000", "000100000", "000100000", "000100000", "000100000",
"000100001", "000100001", "000100001", "000100001", "000100001",
"000100001", "000100010", "000100010", "000100010", "000100010",
"000100010", "000100010", "000100011", "000100011", "000100011",
"000100011", "000100011", "000100011", "000100011", "000100100",
"000100100", "000100100", "000100100", "000100100", "000100100",
"000100101", "000100101", "000100101", "000100101", "000100101",
"000100101", "000100101", "000100110", "000100110", "000100110",
"000100110", "000100110", "000100110", "000100110", "000100111",
"000100111", "000100111", "000100111", "000100111", "000100111",
"000100111", "000101000", "000101000", "000101000", "000101000",
"000101000", "000101000", "000101000", "000101000", "000101001",
"000101001", "000101001", "000101001", "000101001", "000101001",
"000101001", "000101001", "000101010", "000101010", "000101010",
"000101010", "000101010", "000101010", "000101010", "000101010",
"000101011", "000101011", "000101011", "000101011", "000101011",
"000101011", "000101011", "000101011", "000101011", "000101100",
"000101100", "000101100", "000101100", "000101100", "000101100",
"000101100", "000101100", "000101100", "000101101", "000101101",
"000101101", "000101101", "000101101", "000101101", "000101101",
"000101101", "000101101", "000101101", "000101110", "000101110",
"000101110", "000101110", "000101110", "000101110", "000101110",
"000101110", "000101110", "000101110", "000101110", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000101111", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010" );

--table de valeurs pour g�n�rer un sinus de 770 hz
constant sinus770 :defsinus :=( "000000000", "000000001", "000000001", "000000001", "000000001",
"000000010", "000000010", "000000010", "000000010", "000000011",
"000000011", "000000011", "000000011", "000000100", "000000100",
"000000100", "000000100", "000000101", "000000101", "000000101",
"000000101", "000000110", "000000110", "000000110", "000000110",
"000000111", "000000111", "000000111", "000000111", "000000111",
"000001000", "000001000", "000001000", "000001000", "000001001",
"000001001", "000001001", "000001001", "000001010", "000001010",
"000001010", "000001010", "000001011", "000001011", "000001011",
"000001011", "000001100", "000001100", "000001100", "000001100",
"000001100", "000001101", "000001101", "000001101", "000001101",
"000001110", "000001110", "000001110", "000001110", "000001111",
"000001111", "000001111", "000001111", "000010000", "000010000",
"000010000", "000010000", "000010000", "000010001", "000010001",
"000010001", "000010001", "000010010", "000010010", "000010010",
"000010010", "000010010", "000010011", "000010011", "000010011",
"000010011", "000010100", "000010100", "000010100", "000010100",
"000010100", "000010101", "000010101", "000010101", "000010101",
"000010110", "000010110", "000010110", "000010110", "000010110",
"000010111", "000010111", "000010111", "000010111", "000011000",
"000011000", "000011000", "000011000", "000011000", "000011001",
"000011001", "000011001", "000011001", "000011001", "000011010",
"000011010", "000011010", "000011010", "000011010", "000011011",
"000011011", "000011011", "000011011", "000011100", "000011100",
"000011100", "000011100", "000011100", "000011101", "000011101",
"000011101", "000011101", "000011101", "000011110", "000011110",
"000011110", "000011110", "000011110", "000011110", "000011111",
"000011111", "000011111", "000011111", "000011111", "000100000",
"000100000", "000100000", "000100000", "000100000", "000100001",
"000100001", "000100001", "000100001", "000100001", "000100010",
"000100010", "000100010", "000100010", "000100010", "000100010",
"000100011", "000100011", "000100011", "000100011", "000100011",
"000100011", "000100100", "000100100", "000100100", "000100100",
"000100100", "000100100", "000100101", "000100101", "000100101",
"000100101", "000100101", "000100101", "000100110", "000100110",
"000100110", "000100110", "000100110", "000100110", "000100111",
"000100111", "000100111", "000100111", "000100111", "000100111",
"000101000", "000101000", "000101000", "000101000", "000101000",
"000101000", "000101000", "000101001", "000101001", "000101001",
"000101001", "000101001", "000101001", "000101001", "000101010",
"000101010", "000101010", "000101010", "000101010", "000101010",
"000101010", "000101010", "000101011", "000101011", "000101011",
"000101011", "000101011", "000101011", "000101011", "000101100",
"000101100", "000101100", "000101100", "000101100", "000101100",
"000101100", "000101100", "000101100", "000101101", "000101101",
"000101101", "000101101", "000101101", "000101101", "000101101",
"000101101", "000101101", "000101110", "000101110", "000101110",
"000101110", "000101110", "000101110", "000101110", "000101110",
"000101110", "000101110", "000101111", "000101111", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000101111", "000101111", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );

--table de valeurs pour g�n�rer un sinus de 852 hz
constant sinus852 :defsinus :=( "000000000", "000000001", "000000001", "000000001", "000000010",
"000000010", "000000010", "000000010", "000000011", "000000011",
"000000011", "000000011", "000000100", "000000100", "000000100",
"000000101", "000000101", "000000101", "000000101", "000000110",
"000000110", "000000110", "000000110", "000000111", "000000111",
"000000111", "000000111", "000001000", "000001000", "000001000",
"000001000", "000001001", "000001001", "000001001", "000001010",
"000001010", "000001010", "000001010", "000001011", "000001011",
"000001011", "000001011", "000001100", "000001100", "000001100",
"000001100", "000001101", "000001101", "000001101", "000001101",
"000001110", "000001110", "000001110", "000001110", "000001111",
"000001111", "000001111", "000010000", "000010000", "000010000",
"000010000", "000010001", "000010001", "000010001", "000010001",
"000010010", "000010010", "000010010", "000010010", "000010011",
"000010011", "000010011", "000010011", "000010100", "000010100",
"000010100", "000010100", "000010101", "000010101", "000010101",
"000010101", "000010110", "000010110", "000010110", "000010110",
"000010110", "000010111", "000010111", "000010111", "000010111",
"000011000", "000011000", "000011000", "000011000", "000011001",
"000011001", "000011001", "000011001", "000011010", "000011010",
"000011010", "000011010", "000011010", "000011011", "000011011",
"000011011", "000011011", "000011100", "000011100", "000011100",
"000011100", "000011100", "000011101", "000011101", "000011101",
"000011101", "000011110", "000011110", "000011110", "000011110",
"000011110", "000011111", "000011111", "000011111", "000011111",
"000100000", "000100000", "000100000", "000100000", "000100000",
"000100001", "000100001", "000100001", "000100001", "000100001",
"000100010", "000100010", "000100010", "000100010", "000100010",
"000100011", "000100011", "000100011", "000100011", "000100011",
"000100100", "000100100", "000100100", "000100100", "000100100",
"000100100", "000100101", "000100101", "000100101", "000100101",
"000100101", "000100110", "000100110", "000100110", "000100110",
"000100110", "000100110", "000100111", "000100111", "000100111",
"000100111", "000100111", "000100111", "000101000", "000101000",
"000101000", "000101000", "000101000", "000101000", "000101001",
"000101001", "000101001", "000101001", "000101001", "000101001",
"000101010", "000101010", "000101010", "000101010", "000101010",
"000101010", "000101010", "000101011", "000101011", "000101011",
"000101011", "000101011", "000101011", "000101011", "000101100",
"000101100", "000101100", "000101100", "000101100", "000101100",
"000101100", "000101101", "000101101", "000101101", "000101101",
"000101101", "000101101", "000101101", "000101101", "000101101",
"000101110", "000101110", "000101110", "000101110", "000101110",
"000101110", "000101110", "000101110", "000101110", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000101111", "000101111", "000101111", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );

--table de valeurs pour g�n�rer un sinus de 941 hz
constant sinus941 :defsinus :=( "000000000", "000000001", "000000001", "000000001", "000000010",
"000000010", "000000010", "000000011", "000000011", "000000011",
"000000011", "000000100", "000000100", "000000100", "000000101",
"000000101", "000000101", "000000110", "000000110", "000000110",
"000000110", "000000111", "000000111", "000000111", "000001000",
"000001000", "000001000", "000001000", "000001001", "000001001",
"000001001", "000001010", "000001010", "000001010", "000001010",
"000001011", "000001011", "000001011", "000001100", "000001100",
"000001100", "000001101", "000001101", "000001101", "000001101",
"000001110", "000001110", "000001110", "000001111", "000001111",
"000001111", "000001111", "000010000", "000010000", "000010000",
"000010000", "000010001", "000010001", "000010001", "000010010",
"000010010", "000010010", "000010010", "000010011", "000010011",
"000010011", "000010100", "000010100", "000010100", "000010100",
"000010101", "000010101", "000010101", "000010101", "000010110",
"000010110", "000010110", "000010110", "000010111", "000010111",
"000010111", "000011000", "000011000", "000011000", "000011000",
"000011001", "000011001", "000011001", "000011001", "000011010",
"000011010", "000011010", "000011010", "000011011", "000011011",
"000011011", "000011011", "000011100", "000011100", "000011100",
"000011100", "000011101", "000011101", "000011101", "000011101",
"000011110", "000011110", "000011110", "000011110", "000011111",
"000011111", "000011111", "000011111", "000011111", "000100000",
"000100000", "000100000", "000100000", "000100001", "000100001",
"000100001", "000100001", "000100010", "000100010", "000100010",
"000100010", "000100010", "000100011", "000100011", "000100011",
"000100011", "000100011", "000100100", "000100100", "000100100",
"000100100", "000100101", "000100101", "000100101", "000100101",
"000100101", "000100110", "000100110", "000100110", "000100110",
"000100110", "000100110", "000100111", "000100111", "000100111",
"000100111", "000100111", "000101000", "000101000", "000101000",
"000101000", "000101000", "000101001", "000101001", "000101001",
"000101001", "000101001", "000101001", "000101010", "000101010",
"000101010", "000101010", "000101010", "000101010", "000101011",
"000101011", "000101011", "000101011", "000101011", "000101011",
"000101011", "000101100", "000101100", "000101100", "000101100",
"000101100", "000101100", "000101101", "000101101", "000101101",
"000101101", "000101101", "000101101", "000101101", "000101101",
"000101110", "000101110", "000101110", "000101110", "000101110",
"000101110", "000101110", "000101110", "000101111", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000101111", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );

--table de valeurs pour g�n�rer un sinus de 1209 hz
constant sinus1209 :defsinus :=( "000000000", "000000001", "000000001", "000000010", "000000010",
"000000010", "000000011", "000000011", "000000100", "000000100",
"000000100", "000000101", "000000101", "000000101", "000000110",
"000000110", "000000111", "000000111", "000000111", "000001000",
"000001000", "000001000", "000001001", "000001001", "000001010",
"000001010", "000001010", "000001011", "000001011", "000001011",
"000001100", "000001100", "000001101", "000001101", "000001101",
"000001110", "000001110", "000001110", "000001111", "000001111",
"000001111", "000010000", "000010000", "000010001", "000010001",
"000010001", "000010010", "000010010", "000010010", "000010011",
"000010011", "000010011", "000010100", "000010100", "000010100",
"000010101", "000010101", "000010101", "000010110", "000010110",
"000010111", "000010111", "000010111", "000011000", "000011000",
"000011000", "000011001", "000011001", "000011001", "000011010",
"000011010", "000011010", "000011011", "000011011", "000011011",
"000011011", "000011100", "000011100", "000011100", "000011101",
"000011101", "000011101", "000011110", "000011110", "000011110",
"000011111", "000011111", "000011111", "000011111", "000100000",
"000100000", "000100000", "000100001", "000100001", "000100001",
"000100010", "000100010", "000100010", "000100010", "000100011",
"000100011", "000100011", "000100011", "000100100", "000100100",
"000100100", "000100101", "000100101", "000100101", "000100101",
"000100110", "000100110", "000100110", "000100110", "000100111",
"000100111", "000100111", "000100111", "000101000", "000101000",
"000101000", "000101000", "000101000", "000101001", "000101001",
"000101001", "000101001", "000101010", "000101010", "000101010",
"000101010", "000101010", "000101011", "000101011", "000101011",
"000101011", "000101011", "000101100", "000101100", "000101100",
"000101100", "000101100", "000101101", "000101101", "000101101",
"000101101", "000101101", "000101101", "000101110", "000101110",
"000101110", "000101110", "000101110", "000101110", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );

--table de valeurs pour g�n�rer un sinus de 1336 hz
constant sinus1336 : defsinus :=( "000000000", "000000001", "000000001", "000000010", "000000010",
"000000011", "000000011", "000000011", "000000100", "000000100",
"000000101", "000000101", "000000110", "000000110", "000000110",
"000000111", "000000111", "000001000", "000001000", "000001000",
"000001001", "000001001", "000001010", "000001010", "000001011",
"000001011", "000001011", "000001100", "000001100", "000001101",
"000001101", "000001101", "000001110", "000001110", "000001111",
"000001111", "000001111", "000010000", "000010000", "000010001",
"000010001", "000010001", "000010010", "000010010", "000010011",
"000010011", "000010011", "000010100", "000010100", "000010100",
"000010101", "000010101", "000010110", "000010110", "000010110",
"000010111", "000010111", "000011000", "000011000", "000011000",
"000011001", "000011001", "000011001", "000011010", "000011010",
"000011010", "000011011", "000011011", "000011100", "000011100",
"000011100", "000011101", "000011101", "000011101", "000011110",
"000011110", "000011110", "000011111", "000011111", "000011111",
"000100000", "000100000", "000100000", "000100001", "000100001",
"000100001", "000100010", "000100010", "000100010", "000100010",
"000100011", "000100011", "000100011", "000100100", "000100100",
"000100100", "000100101", "000100101", "000100101", "000100101",
"000100110", "000100110", "000100110", "000100111", "000100111",
"000100111", "000100111", "000101000", "000101000", "000101000",
"000101000", "000101001", "000101001", "000101001", "000101001",
"000101010", "000101010", "000101010", "000101010", "000101011",
"000101011", "000101011", "000101011", "000101011", "000101100",
"000101100", "000101100", "000101100", "000101100", "000101101",
"000101101", "000101101", "000101101", "000101101", "000101110",
"000101110", "000101110", "000101110", "000101110", "000101110",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000101111", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );

--table de valeurs pour g�n�rer un sinus de 1477hz
constant sinus1477 :defsinus :=( "000000000", "000000001", "000000001", "000000010", "000000010",
"000000011", "000000011", "000000100", "000000100", "000000101",
"000000101", "000000110", "000000110", "000000111", "000000111",
"000000111", "000001000", "000001000", "000001001", "000001001",
"000001010", "000001010", "000001011", "000001011", "000001100",
"000001100", "000001100", "000001101", "000001101", "000001110",
"000001110", "000001111", "000001111", "000010000", "000010000",
"000010000", "000010001", "000010001", "000010010", "000010010",
"000010011", "000010011", "000010011", "000010100", "000010100",
"000010101", "000010101", "000010110", "000010110", "000010110",
"000010111", "000010111", "000011000", "000011000", "000011001",
"000011001", "000011001", "000011010", "000011010", "000011011",
"000011011", "000011011", "000011100", "000011100", "000011100",
"000011101", "000011101", "000011110", "000011110", "000011110",
"000011111", "000011111", "000011111", "000100000", "000100000",
"000100001", "000100001", "000100001", "000100010", "000100010",
"000100010", "000100011", "000100011", "000100011", "000100100",
"000100100", "000100100", "000100101", "000100101", "000100101",
"000100110", "000100110", "000100110", "000100110", "000100111",
"000100111", "000100111", "000101000", "000101000", "000101000",
"000101001", "000101001", "000101001", "000101001", "000101010",
"000101010", "000101010", "000101010", "000101011", "000101011",
"000101011", "000101011", "000101100", "000101100", "000101100",
"000101100", "000101101", "000101101", "000101101", "000101101",
"000101101", "000101110", "000101110", "000101110", "000101110",
"000101110", "000101111", "000101111", "000101111", "000101111",
"000101111", "000101111", "000110000", "000110000", "000110000",
"000110000", "000110000", "000110000", "000110000", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );

--table de valeurs pour g�n�rer un sinus de 1633 hz
constant sinus1633 :defsinus :=( "000000000", "000000001", "000000010", "000000010", "000000011",
"000000011", "000000100", "000000100", "000000101", "000000101",
"000000110", "000000110", "000000111", "000000111", "000001000",
"000001000", "000001001", "000001001", "000001010", "000001010",
"000001011", "000001011", "000001100", "000001100", "000001101",
"000001101", "000001110", "000001110", "000001111", "000001111",
"000010000", "000010000", "000010001", "000010001", "000010010",
"000010010", "000010011", "000010011", "000010100", "000010100",
"000010100", "000010101", "000010101", "000010110", "000010110",
"000010111", "000010111", "000011000", "000011000", "000011001",
"000011001", "000011001", "000011010", "000011010", "000011011",
"000011011", "000011100", "000011100", "000011101", "000011101",
"000011101", "000011110", "000011110", "000011111", "000011111",
"000011111", "000100000", "000100000", "000100001", "000100001",
"000100001", "000100010", "000100010", "000100011", "000100011",
"000100011", "000100100", "000100100", "000100100", "000100101",
"000100101", "000100101", "000100110", "000100110", "000100110",
"000100111", "000100111", "000100111", "000101000", "000101000",
"000101000", "000101001", "000101001", "000101001", "000101010",
"000101010", "000101010", "000101010", "000101011", "000101011",
"000101011", "000101100", "000101100", "000101100", "000101100",
"000101101", "000101101", "000101101", "000101101", "000101101",
"000101110", "000101110", "000101110", "000101110", "000101111",
"000101111", "000101111", "000101111", "000101111", "000101111",
"000110000", "000110000", "000110000", "000110000", "000110000",
"000110000", "000110001", "000110001", "000110001", "000110001",
"000110001", "000110001", "000110001", "000110001", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000110010", "000110010",
"000110010", "000110010", "000110010", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000", "000000000", "000000000", "000000000",
"000000000", "000000000" );
signal sinus : defsinus;
begin

  -- Process pour sens
  process(rst, h)
    begin
      if(rst='1') then
        sens<='0';
      elsif (h'event and h='1') then
        if C3='1' then sens <= not sens;
        end if;
      end if;
  end process;

  -- Process pour signe
  process(rst, h)
    begin
      if(rst='1') then
        signe<='0';
      elsif (h'event and h='1') then
        if C4='1' then signe <= not signe;
        end if;
      end if;
  end process;

  -- Process pour Vs
  process(rst,h)
      variable mux, mux2 : std_logic_vector(9 downto 0);
       variable flow: defsinus;
       variable fhigh: defsinus ;
  
    begin
      if(rst='1') then
        Vs <=(others => '0');
      elsif (h'event and h='1') then
    case C5 is
      when '0' => mux := 0-('0' & sinusask(conv_integer(I)));
                  mux2 := 0-('0' & sinus(conv_integer(I)));
                  
                  if amp = '0' then
                    mux(8 downto 0) := mux (9 downto 1);
                  end if;
       
      when '1' => mux :=('0' & sinusask(conv_integer(I)));
                  mux2 := ('0' & sinus(conv_integer(I)));
                  
                  if amp = '0' then
                    mux(8 downto 0) := mux (9 downto 1);
                  end if;
        
      when others => mux := (others =>'0');
                     mux2 := (others => '0');
                     
      end case;
      end if;
      
      case mode is 
       when "10" => Vs <= mux;
       when "11" => Vs <= mux2;
       when others => Vs <= "0000000000";
      end case;
  end process;

  -- Process pour I
  process(rst,h)
    begin
      if(rst='1') then
        I<=(others=>'0');
      elsif (h'event and h='1') then
        if C1='1' then I<=I+1;
        elsif C2='1' then I<=I-1;
        end if;
      end if;
  end process;

  process(sens,signe,eq0,eq511)
    begin
      C1<='0';
      C2<='0';
      C3<='0';
      C4<='0';
      C5<='0';
      case std_logic_vector'(sens & signe) is
        when "00" => if eq511='0' then C1<='1';
                                       C5<='1';
                     else C3<='1';
                          C5<='1';
                     end if;
        when "01" => if eq511='0' then C1<='1';
                     else C3<='1';
                     end if;
        when "10" => if eq0='0' then C2<='1';
                                     C5<='1';
                     else C3<='1';
                          C4<='1';
                          C5<='1';
                     end if;
        when others => if eq0='0' then C2<='1';
                       else C3<='1';
                            C4<='1';
                       end if;
      end case;
  end process;

  eq0<='1' when conv_integer(I)=0 else '0';
  eq511<='1' when conv_integer(I)=156 else '0';
  
  
--Processe pour la fr�quence frq
--le d�codage des num�ros se fait dans le contr�leur
--dans le g�n�rateur on positionne juste la bonne fr�quence; ce qui permettra de g�n�rer le bon sinus
--  
process (freq)
  variable flow: defsinus;
  variable fhigh: defsinus ;
  
  begin
    case freq is
  when "0000" => fhigh :=sinus1209;
                 flow  :=sinus697;

  when "0001" => fhigh :=sinus1336;
                 flow :=sinus697;

  when "0010" => fhigh :=sinus1477;
                 flow :=sinus697;

  when "0011" => fhigh :=sinus1633;
                 flow  :=sinus697;

  when "0100" => fhigh :=sinus1209;
                 flow :=sinus770;

  when "0101" => fhigh :=sinus1336;
                 flow :=sinus770;

  when "0110" => fhigh :=sinus1477;
                 flow :=sinus770;

  when "0111" => fhigh :=sinus1633;
                 flow  :=sinus770;

  when "1000" => fhigh :=sinus1209;
                 flow  :=sinus852;

  when "1001" => fhigh :=sinus1336;
                 flow  :=sinus852;

  when "1010" => fhigh :=sinus1477;
                 flow  :=sinus852;

  when "1011" => fhigh :=sinus1633;
                 flow  :=sinus852;

  when "1100" => fhigh :=sinus1209;
                 flow  :=sinus941;

  when "1101" => fhigh :=sinus1336;
                 flow  :=sinus941;

  when "1110" => fhigh :=sinus1477;
                 flow  :=sinus941;

  when "1111" => fhigh :=sinus1633;
                 flow  :=sinus941;
  when others => fhigh :=sinusask;
                 flow  :=sinusask;
  end case;
  
if(fhigh = sinusask ) then sinus <=sinusask;
else 
for i in fhigh'range loop 
  sinus(i) <= std_logic_vector(unsigned(flow(i)) + unsigned(fhigh(i)));
end loop;
end if;
end process;
  
end rtl;

