------------
-- Sine wave ROM
------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity sinus is
  port( rst, h : std_logic;
        Vs : out std_logic_vector(9 downto 0) );
end sinus;

------------
-- ROM architecture
------------

architecture rtl of sinus is

  signal sens, signe, eq511, eq0, C1, C2, C3, C4, C5 : std_logic;
  signal I : std_logic_vector(8 downto 0);
  type defsinus is array(0 to 511) of std_logic_vector(8 downto 0);
  
  constant sinus: defsinus := ("000000000", "000000001", "000000011", "000000100", -- Sine wave ROM
    "000000110","000000111", "000001001", "000001010", "000001100",
    "000001101","000001111", "000010000", "000010010", "000010011",
    "000010101","000010111", "000011000", "000011010", "000011011",
    "000011101","000011110", "000100000", "000100001", "000100011",
    "000100100","000100110", "000100111", "000101001", "000101010",
    "000101100","000101101", "000101111", "000110001", "000110010",
    "000110100","000110101", "000110111", "000111000", "000111010",
    "000111011","000111101", "000111110", "001000000", "001000001",
    "001000011","001000100", "001000110", "001000111", "001001001",
    "001001010","001001100", "001001101", "001001111", "001010000",
    "001010010","001010011", "001010101", "001010110", "001011000",
    "001011010","001011011", "001011101", "001011110", "001100000",
    "001100001","001100011", "001100100", "001100110", "001100111",
    "001101001","001101010", "001101100", "001101101", "001101111",
    "001110000","001110010", "001110011", "001110101", "001110110",
    "001111000","001111001", "001111010", "001111100", "001111101",
    "001111111","010000000", "010000010", "010000011", "010000101",
    "010000110","010001000", "010001001", "010001011", "010001100",
    "010001110","010001111", "010010001", "010010010", "010010100",
    "010010101","010010111", "010011000", "010011001", "010011011",
    "010011100","010011110", "010011111", "010100001", "010100010",
    "010100100","010100101", "010100110", "010101000", "010101001",
    "010101011","010101100", "010101110", "010101111", "010110001",
    "010110010","010110011", "010110101", "010110110", "010111000",
    "010111001","010111011", "010111100", "010111101", "010111111",
    "011000000","011000010", "011000011", "011000100", "011000110",
    "011000111","011001001", "011001010", "011001100", "011001101",
    "011001110","011010000", "011010001", "011010010", "011010100",
    "011010101","011010111", "011011000", "011011001", "011011011",
    "011011100","011011110", "011011111", "011100000", "011100010",
    "011100011","011100100", "011100110", "011100111", "011101000",
    "011101010","011101011", "011101101", "011101110", "011101111",
    "011110001","011110010", "011110011", "011110101", "011110110",
    "011110111","011111001", "011111010", "011111011", "011111101",
    "011111110","011111111", "100000001", "100000010", "100000011",
    "100000100","100000110", "100000111", "100001000", "100001010",
    "100001011","100001100", "100001110", "100001111", "100010000",
    "100010001","100010011", "100010100", "100010101", "100010111",
    "100011000","100011001", "100011010", "100011100", "100011101",
    "100011110","100011111", "100100001", "100100010", "100100011",
    "100100100","100100110", "100100111", "100101000", "100101001",
    "100101011","100101100", "100101101", "100101110", "100101111",
    "100110001","100110010", "100110011", "100110100", "100110110",
    "100110111","100111000", "100111001", "100111010", "100111100",
    "100111101","100111110", "100111111", "101000000", "101000001",
    "101000011","101000100", "101000101", "101000110", "101000111",
    "101001000","101001010", "101001011", "101001100", "101001101",
    "101001110","101001111", "101010000", "101010010", "101010011",
    "101010100","101010101", "101010110", "101010111", "101011000",
    "101011001","101011010", "101011100", "101011101", "101011110",
    "101011111","101100000", "101100001", "101100010", "101100011",
    "101100100","101100101", "101100110", "101101000", "101101001",
    "101101010","101101011", "101101100", "101101101", "101101110",
    "101101111","101110000", "101110001", "101110010", "101110011",
    "101110100","101110101", "101110110", "101110111", "101111000",
    "101111001","101111010", "101111011", "101111100", "101111101",
    "101111110","101111111", "110000000", "110000001", "110000010",
    "110000011","110000100", "110000101", "110000110", "110000111",
    "110001000","110001001", "110001010", "110001011", "110001100",
    "110001100","110001101", "110001110", "110001111", "110010000",
    "110010001","110010010", "110010011", "110010100", "110010101",
    "110010110","110010111", "110010111", "110011000", "110011001",
    "110011010","110011011", "110011100", "110011101", "110011110",
    "110011110","110011111", "110100000", "110100001", "110100010",
    "110100011","110100011", "110100100", "110100101", "110100110",
    "110100111","110101000", "110101000", "110101001", "110101010",
    "110101011","110101100", "110101100", "110101101", "110101110",
    "110101111","110101111", "110110000", "110110001", "110110010",
    "110110011","110110011", "110110100", "110110101", "110110110",
    "110110110","110110111", "110111000", "110111000", "110111001",
    "110111010","110111011", "110111011", "110111100", "110111101",
    "110111101","110111110", "110111111", "110111111", "111000000",
    "111000001","111000010", "111000010", "111000011", "111000011",
    "111000100","111000101", "111000101", "111000110", "111000111",
    "111000111","111001000", "111001001", "111001001", "111001010",
    "111001010","111001011", "111001100", "111001100", "111001101",
    "111001101","111001110", "111001111", "111001111", "111010000",
    "111010000","111010001", "111010001", "111010010", "111010011",
    "111010011","111010100", "111010100", "111010101", "111010101",
    "111010110","111010110", "111010111", "111010111", "111011000",
    "111011000","111011001", "111011001", "111011010", "111011010",
    "111011011","111011011", "111011100", "111011100", "111011101",
    "111011101","111011110", "111011110", "111011110", "111011111",
    "111011111","111100000", "111100000", "111100001", "111100001",
    "111100001","111100010", "111100010", "111100011", "111100011",
    "111100011","111100100", "111100100", "111100101", "111100101",
    "111100101","111100110", "111100110", "111100110", "111100111",
    "111100111","111100111", "111101000", "111101000", "111101000",
    "111101001","111101001", "111101001", "111101010", "111101010",
    "111101010","111101010", "111101011", "111101011", "111101011",
    "111101100","111101100", "111101100", "111101100", "111101101",
    "111101101","111101101", "111101101", "111101110", "111101110",
    "111101110","111101110", "111101111", "111101111", "111101111",
    "111101111","111101111", "111110000", "111110000", "111110000",
    "111110000","111110000", "111110000", "111110001", "111110001",
    "111110001","111110001", "111110001", "111110001", "111110010",
    "111110010","111110010", "111110010", "111110010", "111110010",
    "111110010","111110010", "111110010", "111110011", "111110011",
    "111110011","111110011", "111110011", "111110011", "111110011",
    "111110011","111110011", "111110011", "111110011", "111110011",
    "111110011","111110011", "111110011", "111110011", "111110011",
    "111110011","111110011", "111110011");

  begin

  sens_p: process(rst, h)                      -- Direction process
  begin
    
    if(rst='1') then                           -- On reset
      sens<='0';
    elsif (rising_edge(h)) then                -- On clock rising edge
      if C3='1' then sens <= not sens;         -- Toggle direction on C3
      end if;
    end if;

  end process;

  sign_p: process(rst, h)                      -- Sign process
  begin

    if(rst='1') then                           -- On reset
      signe<='0';
    elsif (rising_edge(h)) then                -- On clock rising edge
      if C4='1' then signe <= not signe;       -- Toggle sign on C4
      end if;
    end if;

  end process;

  vs_p: process(rst, h)                        -- Vs process
  begin

    if(rst='1') then                           -- On reset
      Vs <=(others => '0');
    elsif (rising_edge(h)) then                -- On clock rising edge
      if C5='1' then Vs<=('0' & sinus(conv_integer(I))); -- Output positive waveform on C5, else negative
      else Vs<=0-('0' & sinus(conv_integer(I)));
      end if;
    end if;

  end process;

  i_p: process(rst, h)                         -- Count process
  begin

    if(rst='1') then                           -- On reset
      I<=(others=>'0');
    elsif (rising_edge(h)) then                -- On clock rising edge
      if C1='1' then I<=I+1;                   -- Count up on C1
      elsif C2='1' then I<=I-1;                -- Count down on C2
      end if;
    end if;

  end process;

  state_p: process(sens, signe, eq0, eq511)    -- State process
  begin

    C1<='0';
    C2<='0';
    C3<='0';
    C4<='0';
    C5<='0';

    case std_logic_vector'(sens & signe) is
      when "00" => if eq511='0' then C1<='1';
                                     C5<='1';
                   else C3<='1';
                        C5<='1';
                   end if;
      when "01" => if eq511='0' then C1<='1';
                   else C3<='1';
                   end if;
      when "10" => if eq0='0' then C2<='1';
                                   C5<='1';
                   else C3<='1';
                        C4<='1';
                        C5<='1';
                   end if;
      when others => if eq0='0' then C2<='1';
                     else C3<='1';
                          C4<='1';
                     end if;
    end case;

  end process;

  eq0<='1' when conv_integer(I)=0 else '0';
  eq511<='1' when conv_integer(I)=511 else '0';

end rtl;
