----------------------------------------
----------------------------------------
-------------------
----
--
-- The Von Neumann Calculator
-- A VHDL Project
-- Polytech Nice-Sophia
-- ELEC4
-- 2013
--
----
-------------------
----------------------------------------
----------------------------------------

-- Version 1 : Created the RAM
---- La simulation du RAM a �t� modifi�
---- Au lieu d'utiliser Nbadr = 2**16,
----  nous avons utilis� Nbadr = 2**8
----  car le simulateur n'arrive pas �
----  simuler 63556 case de m�moire

----------------------------------------
------------- Written by ---------------
------ KaiserHaz and Moustapha LO ------
----------------------------------------
----------------------------------------