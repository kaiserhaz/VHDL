----------------------------------------
----------------------------------------
-------------------
----
--
-- RS232 Controller
-- A VHDL Project
-- Polytech Nice-Sophia
-- ELEC5
-- 2013
--
----
-------------------
----------------------------------------
----------------------------------------

entity README is

-- Version 1 : Initially created the RS 232 controller
---- Basically the controller handles RS232 communication
----  with other functionnalities added to it as well

end entity;

----------------------------------------
----------------------------------------
------------- Written by ---------------
----------------------------------------
------------- KaiserHaz ----------------
----------------------------------------
----------------------------------------