----------------------------------------
-- Includes
----------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

----------------------------------------
-- Entite
----------------------------------------

entity sinus is
  port( rst  : in std_logic;
        h    : in std_logic;
        amp  : in std_logic;
        freq : in std_logic_vector(3 downto 0);
        mode : in std_logic_vector(1 downto 0);
        Vs   : out std_logic_vector(9 downto 0) );
end sinus;

----------------------------------------
-- Architecture
----------------------------------------

architecture rtl of sinus is
  
  -- Declaration des signaux
  
  signal sens_ask, sens_dtmf1, sens_dtmf2    : std_logic;
  signal signe_ask, signe_dtmf1, signe_dtmf2 : std_logic;
  signal eqmax_ask, eqmax_dtmf1, eqmax_dtmf2 : std_logic;
  signal supmax_dtmf1, supmax_dtmf2          : std_logic;
  signal eq0_ask, eq0_dtmf1, eq0_dtmf2       : std_logic;
  signal C1_ask, C1_dtmf1, C1_dtmf2          : std_logic;
  signal C2_ask, C2_dtmf1, C2_dtmf2          : std_logic;
  signal C3_ask, C3_dtmf1, C3_dtmf2          : std_logic;
  signal C4_ask, C4_dtmf1, C4_dtmf2          : std_logic;
  signal C5_ask, C5_dtmf1, C5_dtmf2          : std_logic;
  signal C6_ask, C6_dtmf1, C6_dtmf2          : std_logic;
  
  signal I, I1, I2 : integer range 0 to 511 := 0;
  
  signal max1, max2 : integer range 0 to 511 := 0;
  
  signal freq_high, freq_low : std_logic_vector(1 downto 0);
  
  signal tmp_vs : std_logic_vector(9 downto 0);
  
  -- Nouveau type defsinus
 
  type defsinus is array(0 to 357) of std_logic_vector(8 downto 0);
  
  -- Declaration des signaux de type defsinus
  
  signal dtmf_low, dtmf_high : defsinus;
  
  -- Table des valeurs de la porteuse ASK (1600 Hz)
  
  constant sinusask : defsinus :=( "000000000", "000000110", "000001011", "000010000", "000010101",
  "000011010", "000011111", "000100100", "000101001", "000101110",
  "000110011", "000111000", "000111101", "001000010", "001000111",
  "001001100", "001010001", "001010110", "001011010", "001011111",
  "001100100", "001101001", "001101110", "001110011", "001111000",
  "001111101", "010000010", "010000111", "010001011", "010010000",
  "010010101", "010011010", "010011111", "010100011", "010101000",
  "010101101", "010110010", "010110110", "010111011", "011000000",
  "011000100", "011001001", "011001101", "011010010", "011010111",
  "011011011", "011100000", "011100100", "011101001", "011101101",
  "011110001", "011110110", "011111010", "011111110", "100000011",
  "100000111", "100001011", "100010000", "100010100", "100011000",
  "100011100", "100100000", "100100100", "100101000", "100101100",
  "100110000", "100110100", "100111000", "100111100", "101000000",
  "101000100", "101001000", "101001100", "101001111", "101010011",
  "101010111", "101011010", "101011110", "101100010", "101100101",
  "101101001", "101101100", "101110000", "101110011", "101110110",
  "101111010", "101111101", "110000000", "110000011", "110000111",
  "110001010", "110001101", "110010000", "110010011", "110010110",
  "110011001", "110011100", "110011110", "110100001", "110100100",
  "110100111", "110101001", "110101100", "110101111", "110110001",
  "110110100", "110110110", "110111000", "110111011", "110111101",
  "110111111", "111000010", "111000100", "111000110", "111001000",
  "111001010", "111001100", "111001110", "111010000", "111010010",
  "111010100", "111010101", "111010111", "111011001", "111011010",
  "111011100", "111011110", "111011111", "111100000", "111100010",
  "111100011", "111100100", "111100110", "111100111", "111101000",
  "111101001", "111101010", "111101011", "111101100", "111101101",
  "111101110", "111101111", "111101111", "111110000", "111110001",
  "111110001", "111110010", "111110010", "111110011", "111110011",
  "111110100", "111110100", "111110100", "111110100", "111110100",
  "111110100", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
   
  -- Table des valeurs du ton DTMF (697 Hz)
  
  constant sinus697 : defsinus :=("000000000", "000000001", "000000001", "000000001", "000000001",
  "000000010", "000000010", "000000010", "000000010", "000000010",
  "000000011", "000000011", "000000011", "000000011", "000000100",
  "000000100", "000000100", "000000100", "000000100", "000000101",
  "000000101", "000000101", "000000101", "000000110", "000000110",
  "000000110", "000000110", "000000110", "000000111", "000000111",
  "000000111", "000000111", "000000111", "000001000", "000001000",
  "000001000", "000001000", "000001001", "000001001", "000001001",
  "000001001", "000001001", "000001010", "000001010", "000001010",
  "000001010", "000001011", "000001011", "000001011", "000001011",
  "000001011", "000001100", "000001100", "000001100", "000001100",
  "000001100", "000001101", "000001101", "000001101", "000001101",
  "000001101", "000001110", "000001110", "000001110", "000001110",
  "000001111", "000001111", "000001111", "000001111", "000001111",
  "000010000", "000010000", "000010000", "000010000", "000010000",
  "000010001", "000010001", "000010001", "000010001", "000010001",
  "000010010", "000010010", "000010010", "000010010", "000010010",
  "000010011", "000010011", "000010011", "000010011", "000010011",
  "000010100", "000010100", "000010100", "000010100", "000010101",
  "000010101", "000010101", "000010101", "000010101", "000010110",
  "000010110", "000010110", "000010110", "000010110", "000010110",
  "000010111", "000010111", "000010111", "000010111", "000010111",
  "000011000", "000011000", "000011000", "000011000", "000011000",
  "000011001", "000011001", "000011001", "000011001", "000011001",
  "000011010", "000011010", "000011010", "000011010", "000011010",
  "000011011", "000011011", "000011011", "000011011", "000011011",
  "000011011", "000011100", "000011100", "000011100", "000011100",
  "000011100", "000011101", "000011101", "000011101", "000011101",
  "000011101", "000011101", "000011110", "000011110", "000011110",
  "000011110", "000011110", "000011111", "000011111", "000011111",
  "000011111", "000011111", "000011111", "000100000", "000100000",
  "000100000", "000100000", "000100000", "000100000", "000100001",
  "000100001", "000100001", "000100001", "000100001", "000100001",
  "000100010", "000100010", "000100010", "000100010", "000100010",
  "000100010", "000100011", "000100011", "000100011", "000100011",
  "000100011", "000100011", "000100011", "000100100", "000100100",
  "000100100", "000100100", "000100100", "000100100", "000100101",
  "000100101", "000100101", "000100101", "000100101", "000100101",
  "000100101", "000100110", "000100110", "000100110", "000100110",
  "000100110", "000100110", "000100110", "000100111", "000100111",
  "000100111", "000100111", "000100111", "000100111", "000100111",
  "000101000", "000101000", "000101000", "000101000", "000101000",
  "000101000", "000101000", "000101001", "000101001", "000101001",
  "000101001", "000101001", "000101001", "000101001", "000101001",
  "000101010", "000101010", "000101010", "000101010", "000101010",
  "000101010", "000101010", "000101010", "000101011", "000101011",
  "000101011", "000101011", "000101011", "000101011", "000101011",
  "000101011", "000101011", "000101100", "000101100", "000101100",
  "000101100", "000101100", "000101100", "000101100", "000101100",
  "000101100", "000101101", "000101101", "000101101", "000101101",
  "000101101", "000101101", "000101101", "000101101", "000101101",
  "000101101", "000101110", "000101110", "000101110", "000101110",
  "000101110", "000101110", "000101110", "000101110", "000101110",
  "000101110", "000101110", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010" );
  
  -- Table des valeurs du ton DTMF (770 Hz)
  
  constant sinus770 : defsinus :=( "000000000", "000000001", "000000001", "000000001", "000000001",
  "000000010", "000000010", "000000010", "000000010", "000000011",
  "000000011", "000000011", "000000011", "000000100", "000000100",
  "000000100", "000000100", "000000101", "000000101", "000000101",
  "000000101", "000000110", "000000110", "000000110", "000000110",
  "000000111", "000000111", "000000111", "000000111", "000000111",
  "000001000", "000001000", "000001000", "000001000", "000001001",
  "000001001", "000001001", "000001001", "000001010", "000001010",
  "000001010", "000001010", "000001011", "000001011", "000001011",
  "000001011", "000001100", "000001100", "000001100", "000001100",
  "000001100", "000001101", "000001101", "000001101", "000001101",
  "000001110", "000001110", "000001110", "000001110", "000001111",
  "000001111", "000001111", "000001111", "000010000", "000010000",
  "000010000", "000010000", "000010000", "000010001", "000010001",
  "000010001", "000010001", "000010010", "000010010", "000010010",
  "000010010", "000010010", "000010011", "000010011", "000010011",
  "000010011", "000010100", "000010100", "000010100", "000010100",
  "000010100", "000010101", "000010101", "000010101", "000010101",
  "000010110", "000010110", "000010110", "000010110", "000010110",
  "000010111", "000010111", "000010111", "000010111", "000011000",
  "000011000", "000011000", "000011000", "000011000", "000011001",
  "000011001", "000011001", "000011001", "000011001", "000011010",
  "000011010", "000011010", "000011010", "000011010", "000011011",
  "000011011", "000011011", "000011011", "000011100", "000011100",
  "000011100", "000011100", "000011100", "000011101", "000011101",
  "000011101", "000011101", "000011101", "000011110", "000011110",
  "000011110", "000011110", "000011110", "000011110", "000011111",
  "000011111", "000011111", "000011111", "000011111", "000100000",
  "000100000", "000100000", "000100000", "000100000", "000100001",
  "000100001", "000100001", "000100001", "000100001", "000100010",
  "000100010", "000100010", "000100010", "000100010", "000100010",
  "000100011", "000100011", "000100011", "000100011", "000100011",
  "000100011", "000100100", "000100100", "000100100", "000100100",
  "000100100", "000100100", "000100101", "000100101", "000100101",
  "000100101", "000100101", "000100101", "000100110", "000100110",
  "000100110", "000100110", "000100110", "000100110", "000100111",
  "000100111", "000100111", "000100111", "000100111", "000100111",
  "000101000", "000101000", "000101000", "000101000", "000101000",
  "000101000", "000101000", "000101001", "000101001", "000101001",
  "000101001", "000101001", "000101001", "000101001", "000101010",
  "000101010", "000101010", "000101010", "000101010", "000101010",
  "000101010", "000101010", "000101011", "000101011", "000101011",
  "000101011", "000101011", "000101011", "000101011", "000101100",
  "000101100", "000101100", "000101100", "000101100", "000101100",
  "000101100", "000101100", "000101100", "000101101", "000101101",
  "000101101", "000101101", "000101101", "000101101", "000101101",
  "000101101", "000101101", "000101110", "000101110", "000101110",
  "000101110", "000101110", "000101110", "000101110", "000101110",
  "000101110", "000101110", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000101111", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
  -- Table des valeurs du ton DTMF (852 hz)

  constant sinus852 : defsinus :=( "000000000", "000000001", "000000001", "000000001", "000000010",
  "000000010", "000000010", "000000010", "000000011", "000000011",
  "000000011", "000000011", "000000100", "000000100", "000000100",
  "000000101", "000000101", "000000101", "000000101", "000000110",
  "000000110", "000000110", "000000110", "000000111", "000000111",
  "000000111", "000000111", "000001000", "000001000", "000001000",
  "000001000", "000001001", "000001001", "000001001", "000001010",
  "000001010", "000001010", "000001010", "000001011", "000001011",
  "000001011", "000001011", "000001100", "000001100", "000001100",
  "000001100", "000001101", "000001101", "000001101", "000001101",
  "000001110", "000001110", "000001110", "000001110", "000001111",
  "000001111", "000001111", "000010000", "000010000", "000010000",
  "000010000", "000010001", "000010001", "000010001", "000010001",
  "000010010", "000010010", "000010010", "000010010", "000010011",
  "000010011", "000010011", "000010011", "000010100", "000010100",
  "000010100", "000010100", "000010101", "000010101", "000010101",
  "000010101", "000010110", "000010110", "000010110", "000010110",
  "000010110", "000010111", "000010111", "000010111", "000010111",
  "000011000", "000011000", "000011000", "000011000", "000011001",
  "000011001", "000011001", "000011001", "000011010", "000011010",
  "000011010", "000011010", "000011010", "000011011", "000011011",
  "000011011", "000011011", "000011100", "000011100", "000011100",
  "000011100", "000011100", "000011101", "000011101", "000011101",
  "000011101", "000011110", "000011110", "000011110", "000011110",
  "000011110", "000011111", "000011111", "000011111", "000011111",
  "000100000", "000100000", "000100000", "000100000", "000100000",
  "000100001", "000100001", "000100001", "000100001", "000100001",
  "000100010", "000100010", "000100010", "000100010", "000100010",
  "000100011", "000100011", "000100011", "000100011", "000100011",
  "000100100", "000100100", "000100100", "000100100", "000100100",
  "000100100", "000100101", "000100101", "000100101", "000100101",
  "000100101", "000100110", "000100110", "000100110", "000100110",
  "000100110", "000100110", "000100111", "000100111", "000100111",
  "000100111", "000100111", "000100111", "000101000", "000101000",
  "000101000", "000101000", "000101000", "000101000", "000101001",
  "000101001", "000101001", "000101001", "000101001", "000101001",
  "000101010", "000101010", "000101010", "000101010", "000101010",
  "000101010", "000101010", "000101011", "000101011", "000101011",
  "000101011", "000101011", "000101011", "000101011", "000101100",
  "000101100", "000101100", "000101100", "000101100", "000101100",
  "000101100", "000101101", "000101101", "000101101", "000101101",
  "000101101", "000101101", "000101101", "000101101", "000101101",
  "000101110", "000101110", "000101110", "000101110", "000101110",
  "000101110", "000101110", "000101110", "000101110", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
  -- Table des valeurs du ton DTMF (941 Hz)
  
  constant sinus941 : defsinus :=("000000000", "000000001", "000000001", "000000001", "000000010",
  "000000010", "000000010", "000000011", "000000011", "000000011",
  "000000011", "000000100", "000000100", "000000100", "000000101",
  "000000101", "000000101", "000000110", "000000110", "000000110",
  "000000110", "000000111", "000000111", "000000111", "000001000",
  "000001000", "000001000", "000001000", "000001001", "000001001",
  "000001001", "000001010", "000001010", "000001010", "000001010",
  "000001011", "000001011", "000001011", "000001100", "000001100",
  "000001100", "000001101", "000001101", "000001101", "000001101",
  "000001110", "000001110", "000001110", "000001111", "000001111",
  "000001111", "000001111", "000010000", "000010000", "000010000",
  "000010000", "000010001", "000010001", "000010001", "000010010",
  "000010010", "000010010", "000010010", "000010011", "000010011",
  "000010011", "000010100", "000010100", "000010100", "000010100",
  "000010101", "000010101", "000010101", "000010101", "000010110",
  "000010110", "000010110", "000010110", "000010111", "000010111",
  "000010111", "000011000", "000011000", "000011000", "000011000",
  "000011001", "000011001", "000011001", "000011001", "000011010",
  "000011010", "000011010", "000011010", "000011011", "000011011",
  "000011011", "000011011", "000011100", "000011100", "000011100",
  "000011100", "000011101", "000011101", "000011101", "000011101",
  "000011110", "000011110", "000011110", "000011110", "000011111",
  "000011111", "000011111", "000011111", "000011111", "000100000",
  "000100000", "000100000", "000100000", "000100001", "000100001",
  "000100001", "000100001", "000100010", "000100010", "000100010",
  "000100010", "000100010", "000100011", "000100011", "000100011",
  "000100011", "000100011", "000100100", "000100100", "000100100",
  "000100100", "000100101", "000100101", "000100101", "000100101",
  "000100101", "000100110", "000100110", "000100110", "000100110",
  "000100110", "000100110", "000100111", "000100111", "000100111",
  "000100111", "000100111", "000101000", "000101000", "000101000",
  "000101000", "000101000", "000101001", "000101001", "000101001",
  "000101001", "000101001", "000101001", "000101010", "000101010",
  "000101010", "000101010", "000101010", "000101010", "000101011",
  "000101011", "000101011", "000101011", "000101011", "000101011",
  "000101011", "000101100", "000101100", "000101100", "000101100",
  "000101100", "000101100", "000101101", "000101101", "000101101",
  "000101101", "000101101", "000101101", "000101101", "000101101",
  "000101110", "000101110", "000101110", "000101110", "000101110",
  "000101110", "000101110", "000101110", "000101111", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
  -- Table des valeurs du ton DTMF (1209 Hz)
  
  constant sinus1209 : defsinus :=("000000000", "000000001", "000000001", "000000010", "000000010",
  "000000010", "000000011", "000000011", "000000100", "000000100",
  "000000100", "000000101", "000000101", "000000101", "000000110",
  "000000110", "000000111", "000000111", "000000111", "000001000",
  "000001000", "000001000", "000001001", "000001001", "000001010",
  "000001010", "000001010", "000001011", "000001011", "000001011",
  "000001100", "000001100", "000001101", "000001101", "000001101",
  "000001110", "000001110", "000001110", "000001111", "000001111",
  "000001111", "000010000", "000010000", "000010001", "000010001",
  "000010001", "000010010", "000010010", "000010010", "000010011",
  "000010011", "000010011", "000010100", "000010100", "000010100",
  "000010101", "000010101", "000010101", "000010110", "000010110",
  "000010111", "000010111", "000010111", "000011000", "000011000",
  "000011000", "000011001", "000011001", "000011001", "000011010",
  "000011010", "000011010", "000011011", "000011011", "000011011",
  "000011011", "000011100", "000011100", "000011100", "000011101",
  "000011101", "000011101", "000011110", "000011110", "000011110",
  "000011111", "000011111", "000011111", "000011111", "000100000",
  "000100000", "000100000", "000100001", "000100001", "000100001",
  "000100010", "000100010", "000100010", "000100010", "000100011",
  "000100011", "000100011", "000100011", "000100100", "000100100",
  "000100100", "000100101", "000100101", "000100101", "000100101",
  "000100110", "000100110", "000100110", "000100110", "000100111",
  "000100111", "000100111", "000100111", "000101000", "000101000",
  "000101000", "000101000", "000101000", "000101001", "000101001",
  "000101001", "000101001", "000101010", "000101010", "000101010",
  "000101010", "000101010", "000101011", "000101011", "000101011",
  "000101011", "000101011", "000101100", "000101100", "000101100",
  "000101100", "000101100", "000101101", "000101101", "000101101",
  "000101101", "000101101", "000101101", "000101110", "000101110",
  "000101110", "000101110", "000101110", "000101110", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
  -- Table des valeurs du ton DTMF (1336 Hz)
  
  constant sinus1336 : defsinus := ( "000000000", "000000001", "000000001", "000000010", "000000010",
  "000000011", "000000011", "000000011", "000000100", "000000100",
  "000000101", "000000101", "000000110", "000000110", "000000110",
  "000000111", "000000111", "000001000", "000001000", "000001000",
  "000001001", "000001001", "000001010", "000001010", "000001011",
  "000001011", "000001011", "000001100", "000001100", "000001101",
  "000001101", "000001101", "000001110", "000001110", "000001111",
  "000001111", "000001111", "000010000", "000010000", "000010001",
  "000010001", "000010001", "000010010", "000010010", "000010011",
  "000010011", "000010011", "000010100", "000010100", "000010100",
  "000010101", "000010101", "000010110", "000010110", "000010110",
  "000010111", "000010111", "000011000", "000011000", "000011000",
  "000011001", "000011001", "000011001", "000011010", "000011010",
  "000011010", "000011011", "000011011", "000011100", "000011100",
  "000011100", "000011101", "000011101", "000011101", "000011110",
  "000011110", "000011110", "000011111", "000011111", "000011111",
  "000100000", "000100000", "000100000", "000100001", "000100001",
  "000100001", "000100010", "000100010", "000100010", "000100010",
  "000100011", "000100011", "000100011", "000100100", "000100100",
  "000100100", "000100101", "000100101", "000100101", "000100101",
  "000100110", "000100110", "000100110", "000100111", "000100111",
  "000100111", "000100111", "000101000", "000101000", "000101000",
  "000101000", "000101001", "000101001", "000101001", "000101001",
  "000101010", "000101010", "000101010", "000101010", "000101011",
  "000101011", "000101011", "000101011", "000101011", "000101100",
  "000101100", "000101100", "000101100", "000101100", "000101101",
  "000101101", "000101101", "000101101", "000101101", "000101110",
  "000101110", "000101110", "000101110", "000101110", "000101110",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
  -- Table des valeurs du ton DTMF (1477 Hz)
  
  constant sinus1477 : defsinus :=("000000000", "000000001", "000000001", "000000010", "000000010",
  "000000011", "000000011", "000000100", "000000100", "000000101",
  "000000101", "000000110", "000000110", "000000111", "000000111",
  "000000111", "000001000", "000001000", "000001001", "000001001",
  "000001010", "000001010", "000001011", "000001011", "000001100",
  "000001100", "000001100", "000001101", "000001101", "000001110",
  "000001110", "000001111", "000001111", "000010000", "000010000",
  "000010000", "000010001", "000010001", "000010010", "000010010",
  "000010011", "000010011", "000010011", "000010100", "000010100",
  "000010101", "000010101", "000010110", "000010110", "000010110",
  "000010111", "000010111", "000011000", "000011000", "000011001",
  "000011001", "000011001", "000011010", "000011010", "000011011",
  "000011011", "000011011", "000011100", "000011100", "000011100",
  "000011101", "000011101", "000011110", "000011110", "000011110",
  "000011111", "000011111", "000011111", "000100000", "000100000",
  "000100001", "000100001", "000100001", "000100010", "000100010",
  "000100010", "000100011", "000100011", "000100011", "000100100",
  "000100100", "000100100", "000100101", "000100101", "000100101",
  "000100110", "000100110", "000100110", "000100110", "000100111",
  "000100111", "000100111", "000101000", "000101000", "000101000",
  "000101001", "000101001", "000101001", "000101001", "000101010",
  "000101010", "000101010", "000101010", "000101011", "000101011",
  "000101011", "000101011", "000101100", "000101100", "000101100",
  "000101100", "000101101", "000101101", "000101101", "000101101",
  "000101101", "000101110", "000101110", "000101110", "000101110",
  "000101110", "000101111", "000101111", "000101111", "000101111",
  "000101111", "000101111", "000110000", "000110000", "000110000",
  "000110000", "000110000", "000110000", "000110000", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
  -- Table des valeurs du ton DTMF (1633 Hz)
  
  constant sinus1633 :defsinus :=( "000000000", "000000001", "000000010", "000000010", "000000011",
  "000000011", "000000100", "000000100", "000000101", "000000101",
  "000000110", "000000110", "000000111", "000000111", "000001000",
  "000001000", "000001001", "000001001", "000001010", "000001010",
  "000001011", "000001011", "000001100", "000001100", "000001101",
  "000001101", "000001110", "000001110", "000001111", "000001111",
  "000010000", "000010000", "000010001", "000010001", "000010010",
  "000010010", "000010011", "000010011", "000010100", "000010100",
  "000010100", "000010101", "000010101", "000010110", "000010110",
  "000010111", "000010111", "000011000", "000011000", "000011001",
  "000011001", "000011001", "000011010", "000011010", "000011011",
  "000011011", "000011100", "000011100", "000011101", "000011101",
  "000011101", "000011110", "000011110", "000011111", "000011111",
  "000011111", "000100000", "000100000", "000100001", "000100001",
  "000100001", "000100010", "000100010", "000100011", "000100011",
  "000100011", "000100100", "000100100", "000100100", "000100101",
  "000100101", "000100101", "000100110", "000100110", "000100110",
  "000100111", "000100111", "000100111", "000101000", "000101000",
  "000101000", "000101001", "000101001", "000101001", "000101010",
  "000101010", "000101010", "000101010", "000101011", "000101011",
  "000101011", "000101100", "000101100", "000101100", "000101100",
  "000101101", "000101101", "000101101", "000101101", "000101101",
  "000101110", "000101110", "000101110", "000101110", "000101111",
  "000101111", "000101111", "000101111", "000101111", "000101111",
  "000110000", "000110000", "000110000", "000110000", "000110000",
  "000110000", "000110001", "000110001", "000110001", "000110001",
  "000110001", "000110001", "000110001", "000110001", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000110010", "000110010",
  "000110010", "000110010", "000110010", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000", "000000000", "000000000",
  "000000000", "000000000", "000000000" );
  
begin

  ----------------------------------------
  -- Process pour sens
  ----------------------------------------
  
  --- ASK
  
  sens_ask_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      sens_ask <= '0';
      
    elsif (h'event and h='1') then
      if(C3_ask='1') then
        sens_ask <= not sens_ask;
      
      end if;
      
    end if;
    
  end process;
  
  --- DTMF1
  
  sens_dtmf1_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      sens_dtmf1 <= '0';
      
    elsif (h'event and h='1') then
      if(C3_dtmf1='1') then
        sens_dtmf1 <= not sens_dtmf1;
        
      end if;
      
    end if;
    
  end process;
  
  --- DTMF2
  
  sens_dtmf2_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      sens_dtmf2 <= '0';
      
    elsif (h'event and h='1') then       
      if(C3_dtmf2='1') then
        sens_dtmf2 <= not sens_dtmf2;
        
      end if;
      
    end if;
    
  end process;

  ----------------------------------------
  -- Process pour signe
  ----------------------------------------
  
  --- ASK
  
  signe_ask_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      signe_ask <= '0';
      
    elsif (h'event and h='1') then
      if(C4_ask='1') then
        signe_ask <= not signe_ask;
        
      end if;
      
    end if;
    
  end process;
  
  --- DTMF1
  
  signe_dtmf1_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      signe_dtmf1 <= '0';
      
    elsif (h'event and h='1') then
      if(C4_dtmf1='1') then
        signe_dtmf1 <= not signe_dtmf1;
        
      end if;
      
    end if;
    
  end process;
  
  --- DTMF2
  
  signe_dtmf2_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      signe_dtmf2 <= '0';
      
    elsif (h'event and h='1') then      
      if(C4_dtmf2='1') then
        signe_dtmf2 <= not signe_dtmf2;
        
      end if;
      
    end if;
    
  end process;

  ----------------------------------------
  -- Process pour Vs
  ----------------------------------------
  
  vs_p:process(rst, h)
    
    variable mux, mux2 : std_logic_vector(9 downto 0) := "0000000000";
  
  begin
    
    if(rst='1') then
      mux := (others => '0');
      mux2 := (others => '0');
      
    elsif (h'event and h='1') then      
      if(C6_ask = '0') then
        mux := ('0' & sinusask(I));
      
        case C5_ask is
          when '0' => mux := 0 - mux;
          when '1' => mux := mux;
          when others => mux := (others =>'0');
                       
        end case;
        
        if amp = '0' then
          mux(8 downto 0) := mux (9 downto 1);
        end if;
        
        tmp_vs <= mux;
        
      elsif(C6_dtmf1='0' and C6_dtmf2='0') then
        mux := ('0' & dtmf_high(I1));
        mux2 := ('0' & dtmf_low(I2));
      
        case C5_dtmf1 is
          when '0' => mux := 0 - mux;
          when '1' => mux := mux;
          when others => mux := (others =>'0');
                       
        end case;
        
        case C5_dtmf2 is
          when '0' => mux2 := 0 - mux2;         
          when '1' => mux2 := mux2;
          when others => mux2 := (others => '0');
                       
        end case;
        
        tmp_vs <= mux +  mux2;
        
      else
        mux := (others => '0');
        mux2 := (others => '0');
        
        tmp_vs <= (others => '0');
        
      end if;
      
    end if;
          
  end process;

  ----------------------------------------
  -- Process pour I
  ----------------------------------------
  
  i_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      I <= 0;
      
    elsif (h'event and h='1') then
      if(C6_ask='1') then
        I <= 0;
        
      elsif(C1_ask='1') then
        I <= I+1;
        
      elsif(C2_ask='1') then
        I <= I-1;
        
      end if;
      
    end if;
    
  end process;
  
  ----------------------------------------
  -- Process pour I1
  ----------------------------------------
  
  i1_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      I1 <= 0;
      
    elsif (h'event and h='1') then
      if(C6_dtmf1='1') then
        I1 <= 0;
        
      elsif(C1_dtmf1='1') then
        I1 <= I1+1;
        
      elsif(C2_dtmf1='1') then
        I1 <= I1-1;
        
      end if;
      
    end if;
    
  end process;
  
  ----------------------------------------
  -- Process pour I2
  ----------------------------------------
  
  i2_p:process(rst, h)
    
  begin
    
    if(rst='1') then
      I2 <= 0;
      
    elsif (h'event and h='1') then
      if(C6_dtmf2='1') then
        I2 <= 0;
        
      elsif(C1_dtmf2='1') then
        I2 <= I2+1;
        
      elsif(C2_dtmf2='1') then
        I2 <= I2-1;
        
      end if;
      
    end if;
    
  end process;

  ----------------------------------------
  -- Process pour signaux de controles
  ----------------------------------------

  --- ASK

  sig_ask_p:process(sens_ask, signe_ask, eq0_ask, eqmax_ask)
    
    variable ss : std_logic_vector(1 downto 0);
    
  begin
    
    C1_ask <= '0';
    C2_ask <= '0';
    C3_ask <= '0';
    C4_ask <= '0';
    C5_ask <= '0';
    
    ss := sens_ask & signe_ask;

    case ss is
      when "00" => if eqmax_ask='0' then
                    C1_ask<='1';
                    C5_ask<='1';
                    
                   else
                    C3_ask<='1';
                    C5_ask<='1';
                    
                   end if;
                   
      when "01" => if eqmax_ask='0' then
                    C1_ask<='1';
                    
                   else
                    C3_ask<='1';
                    
                   end if;
                   
      when "10" => if eq0_ask='0' then
                    C2_ask<='1';
                    C5_ask<='1';
                    
                   else
                    C3_ask<='1';
                    C4_ask<='1';
                    C5_ask<='1';
                    
                   end if;
                   
      when others => if eq0_ask='0' then
                      C2_ask<='1';
                      
                     else
                      C3_ask<='1';
                      C4_ask<='1';
                      
                     end if;
                     
    end case;
    
  end process;
  
  -- DTMF1

  sig_dtmf1_p:process(sens_dtmf1, signe_dtmf1, eq0_dtmf1, eqmax_dtmf1, supmax_dtmf1)
    
    variable ss : std_logic_vector(1 downto 0);
    
  begin
    
    C1_dtmf1 <= '0';
    C2_dtmf1 <= '0';
    C3_dtmf1 <= '0';
    C4_dtmf1 <= '0';
    C5_dtmf1 <= '0';
    C6_dtmf1 <= '0';
    
    ss := sens_dtmf1 & signe_dtmf1;
    
    if(supmax_dtmf1='1') then
      C6_dtmf1 <= '1';
    
    end if;

    case ss is
      when "00" => if eqmax_dtmf1='0' then
                    C1_dtmf1<='1';
                    C5_dtmf1<='1';
                    
                   else
                    C3_dtmf1<='1';
                    C5_dtmf1<='1';
                    
                   end if;
                   
      when "01" => if eqmax_dtmf1='0' then
                    C1_dtmf1<='1';
                    
                   else
                    C3_dtmf1<='1';
                    
                   end if;
                   
      when "10" => if eq0_dtmf1='0' then
                    C2_dtmf1<='1';
                    C5_dtmf1<='1';
                    
                   else
                    C3_dtmf1<='1';
                    C4_dtmf1<='1';
                    C5_dtmf1<='1';
                    
                   end if;
                   
      when others => if eq0_dtmf1='0' then
                      C2_dtmf1<='1';
                      
                     else
                      C3_dtmf1<='1';
                      C4_dtmf1<='1';
                      
                     end if;
                     
    end case;

  end process;
  
  -- DTMF2

  sig_dtmf2_p:process(sens_dtmf2, signe_dtmf2, eq0_dtmf2, eqmax_dtmf2, supmax_dtmf2)
    
    variable ss : std_logic_vector(1 downto 0);
    
  begin
    
    C1_dtmf2 <= '0';
    C2_dtmf2 <= '0';
    C3_dtmf2 <= '0';
    C4_dtmf2 <= '0';
    C5_dtmf2 <= '0';
    C6_dtmf2 <= '0';
    
    ss := sens_dtmf2 & signe_dtmf2;
    
    if(supmax_dtmf2='1') then
      C6_dtmf2 <= '1';
    
    end if;
    
    case ss is
      when "00" => if eqmax_dtmf2='0' then
                    C1_dtmf2<='1';
                    C5_dtmf2<='1';
                    
                   else
                    C3_dtmf2<='1';
                    C5_dtmf2<='1';
                    
                   end if;
                   
      when "01" => if eqmax_dtmf2='0' then
                    C1_dtmf2<='1';
                    
                   else
                    C3_dtmf2<='1';
                    
                   end if;
                   
      when "10" => if eq0_dtmf2='0' then
                    C2_dtmf2<='1';
                    C5_dtmf2<='1';
                    
                   else
                    C3_dtmf2<='1';
                    C4_dtmf2<='1';
                    C5_dtmf2<='1';
                    
                   end if;
                   
      when others => if eq0_dtmf2='0' then
                      C2_dtmf2<='1';
                      
                     else
                      C3_dtmf2<='1';
                      C4_dtmf2<='1';
                      
                     end if;
                     
    end case;

  end process;
  
  ----------------------------------------
  -- Process pour mode
  ----------------------------------------
  
  mode_p:process(mode)
  
  begin
    
    case mode(0) is
      
      when '0' => C6_ask <= '0';
                  
      when '1' => C6_ask <= '1';
                  
      when others => C6_ask <= '0';
                     
    end case;
    
  end process;
  
  ----------------------------------------
  -- Process pour freq
  ----------------------------------------
  
  freq_p:process(freq)
  
  begin
    
    case freq is
      
    when "0000" => freq_high <= "00";
                   freq_low <= "00";
                   
    when "0001" => freq_high <= "00";
                   freq_low <= "01";
    
    when "0010" => freq_high <= "00";
                   freq_low <= "10";
    
    when "0011" => freq_high <= "00";
                   freq_low <= "11";
    
    when "0100" => freq_high <= "01";
                   freq_low <= "00";
    
    when "0101" => freq_high <= "01";
                   freq_low <= "01";
                   
    when "0110" => freq_high <= "01";
                   freq_low <= "10";
                   
    when "0111" => freq_high <= "01";
                   freq_low <= "11";
                   
    when "1000" => freq_high <= "10";
                   freq_low <= "00";
                   
    when "1001" => freq_high <= "10";
                   freq_low <= "01";
                   
    when "1010" => freq_high <= "10";
                   freq_low <= "10";
                   
    when "1011" => freq_high <= "10";
                   freq_low <= "11";
    
    when "1100" => freq_high <= "11";
                   freq_low <= "00";
                   
    when "1101" => freq_high <= "11";
                   freq_low <= "01";
                   
    when "1110" => freq_high <= "11";
                   freq_low <= "10";
                   
    when "1111" => freq_high <= "11";
                   freq_low <= "11";
                   
    when others => freq_high <= "00";
                   freq_low <= "00";
                   
    end case;
    
  end process;
  
  ----------------------------------------
  -- Process pour dtmf_high
  ----------------------------------------
   
  dtmf_high_p:process(freq_high)
  
  begin
    
    case freq_high is
      
      when "00" => dtmf_high <= sinus1209;
      when "01" => dtmf_high <= sinus1336;
      when "10" => dtmf_high <= sinus1477;
      when "11" => dtmf_high <= sinus1633;
      when others => dtmf_high <= sinus1209;
        
    end case;
    
  end process;
  
  ----------------------------------------
  -- Process pour dtmf_low
  ----------------------------------------
   
  freq_low_p:process(freq_low)
    
  begin
    
    case freq_low is
      
      when "00" => dtmf_low  <= sinus697;
      when "01" => dtmf_low  <= sinus770;
      when "10" => dtmf_low  <= sinus852;
      when "11" => dtmf_low  <= sinus941;
      when others => dtmf_low  <= sinus697;
                     
    end case;
    
  end process;
  
  ----------------------------------------
  -- Process pour max1
  ----------------------------------------
   
  max_1_p:process(freq_high)
    
  begin
    
    case freq_high is
      
      when "00" => max1 <= 206;
      when "01" => max1 <= 186;
      when "10" => max1 <= 168;
      when "11" => max1 <= 152;
      when others => max1 <= 206;

    end case;
    
  end process;
  
  ----------------------------------------
  -- Process pour max2
  ----------------------------------------
   
  max_2_p:process(freq_low)
    
  begin
    
    case freq_low is
      
      when "00" => max2 <= 357;  
      when "01" => max2 <= 324; 
      when "10" => max2 <= 293;   
      when "11" => max2 <= 265;
      when others => max2 <= 357;
                     
    end case;
    
  end process;
  
  ----------------------------------------
  -- Affectation concurrente
  ----------------------------------------

  eq0_ask <= '1' when I=0 else '0';
  eq0_dtmf1 <= '1' when I1=0 else '0';
  eq0_dtmf2 <= '1' when I2=0 else '0';
  
  eqmax_ask <= '1' when I>=155 else '0';
  eqmax_dtmf1 <= '1' when I1=max1 else '0';
  eqmax_dtmf2 <= '1' when I2=max2 else '0';
  
  supmax_dtmf1 <= '1' when I1>max1 else '0';
  supmax_dtmf2 <= '1' when I2>max2 else '0';
  
  Vs <= tmp_vs when (mode(1)='1') else (others => '0');
  
end rtl;